-- megafunction wizard: %LPM_MULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mult 

-- ============================================================
-- File Name: multiplicacao.vhd
-- Megafunction Name(s):
-- 			lpm_mult
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY multiplicacao IS
	PORT(	dataa		: IN STD_LOGIC_VECTOR (2 DOWNTO 0); 		-- entrada a
			datab		: IN STD_LOGIC_VECTOR (2 DOWNTO 0); 		-- entrada b
			result		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0));	-- resultado
END multiplicacao;

ARCHITECTURE SYN OF multiplicacao IS
-- sinal que é que recebe o resultado do componente lpm_mult
SIGNAL sub_wire0	: STD_LOGIC_VECTOR (5 DOWNTO 0);
-- MEGAFUNCTION: multiplicação
COMPONENT lpm_mult
GENERIC (lpm_hint					: STRING;
			lpm_representation	: STRING;
			lpm_type					: STRING;
			lpm_widtha			: NATURAL;
			lpm_widthb			: NATURAL;
			lpm_widthp			: NATURAL);
	PORT (dataa		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			datab		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (5 DOWNTO 0));
END COMPONENT;

BEGIN
-- atribui o resultado contido no sub_wire0 para o outpu
	result    <= sub_wire0(5 DOWNTO 0);
-- MEGAFUNCTION: multiplicação
	lpm_mult_component : lpm_mult
	GENERIC MAP (
		lpm_hint => "MAXIMIZE_SPEED=5",
		lpm_representation => "UNSIGNED",
		lpm_type => "LPM_MULT",
		lpm_widtha => 3,	-- nº bits de a 
		lpm_widthb => 3,	-- nº bits de b
		lpm_widthp => 6) 	-- largura total 
	PORT MAP ( 	dataa => dataa,			-- a
 					datab => datab,			-- b
					result => sub_wire0); 	-- resultado

END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
-- Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantB NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: SignedMult NUMERIC "0"
-- Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
-- Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
-- Retrieval info: PRIVATE: WidthA NUMERIC "3"
-- Retrieval info: PRIVATE: WidthB NUMERIC "3"
-- Retrieval info: PRIVATE: WidthP NUMERIC "6"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: PRIVATE: optimize NUMERIC "0"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=5"
-- Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
-- Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "3"
-- Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "3"
-- Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "6"
-- Retrieval info: USED_PORT: dataa 0 0 3 0 INPUT NODEFVAL "dataa[2..0]"
-- Retrieval info: USED_PORT: datab 0 0 3 0 INPUT NODEFVAL "datab[2..0]"
-- Retrieval info: USED_PORT: result 0 0 6 0 OUTPUT NODEFVAL "result[5..0]"
-- Retrieval info: CONNECT: @dataa 0 0 3 0 dataa 0 0 3 0
-- Retrieval info: CONNECT: @datab 0 0 3 0 datab 0 0 3 0
-- Retrieval info: CONNECT: result 0 0 6 0 @result 0 0 6 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL multiplicacao.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL multiplicacao.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL multiplicacao.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL multiplicacao.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL multiplicacao_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
